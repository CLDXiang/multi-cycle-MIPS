`timescale 1ns / 1ps

module top(
        input logic clk, reset
    );
endmodule
